///////////////////////////////////////////////////////////////////////////////
// File:        algn_types.sv
// Author:      Ahmed Awad-Allah Mohamed
// Date:        2025-10-12
// Description: Type Definitions for the Alignment Controller Verification Environment
//
// -----------------------------------------------------------------------------
// Overview:
// This file defines common types and aliases used throughout the verification
// environment of the Alignment Controller (ALGN). These definitions serve as 
// shared building blocks between testbench components (e.g., environment, agent,
// monitor, model, and scoreboard).
//
// -----------------------------------------------------------------------------
// Code Flow & Purpose:
// 1. **Virtual Interface Definition**
//    - Declares a `typedef` for the virtual interface `algn_vif`.
//    - This allows any UVM component (e.g., driver, monitor, model) to access 
//      the DUT interface through a consistent handle without hardcoding 
//      the interface type name.
//    - Example usage:
//         algn_vif vif;
//         vif = my_config.get_vif(); // Retrieved via UVM configuration DB.
//
// 2. **IRQ Structure Definition**
//    - Defines a small structure `irq` to represent interrupt-related information
//      observed or generated by the DUT.
//    - It contains:
//         * `irq_value`: logic level of the IRQ line (1 = asserted, 0 = deasserted)
//         * `irq_type`: textual identifier describing the IRQ cause/type 
//                      (e.g., "rx_done", "tx_done", "alignment_error").
//
// 3. **Usage in Environment**
//    - These types are included (via `include "algn_types.sv"`) in multiple 
//      components such as the environment, monitor, or model to ensure type 
//      consistency across the testbench.
//    - The virtual interface handle (`algn_vif`) allows dynamic binding to 
//      different interface instances during simulation setup.
//    - The `irq` struct provides a convenient way to pass interrupt information 
//      between analysis components (monitor → scoreboard/model).
//
// -----------------------------------------------------------------------------
// This file should be included early in the testbench hierarchy (e.g. in env.sv)
// to ensure all components have access to the shared type definitions.
// -----------------------------------------------------------------------------
///////////////////////////////////////////////////////////////////////////////

`ifndef ALGN_TYPES
  `define ALGN_TYPES

  //--------------------------------------------------------------------------
  // Virtual Interface Type
  //--------------------------------------------------------------------------
  // 'algn_vif' is a shorthand alias for the virtual interface of type 'algn_if'.
  // It enables UVM components to connect to the DUT interface through configuration.
  typedef virtual algn_if algn_vif;


  //--------------------------------------------------------------------------
  // IRQ Structure
  //--------------------------------------------------------------------------
  // Represents the state and classification of an interrupt event.
  typedef struct {
    bit     irq_value;   // Actual logic value of the IRQ signal (1 = asserted)
    string  irq_type;    // Descriptive type of the interrupt (e.g., "rx_done")
  } irq;

`endif
