///////////////////////////////////////////////////////////////////////////////
// File:        algn_coverage.sv
// Author:      Ahmed Awad-Allah Mohamed
// Date:        12/10/2025
// Description: Functional Coverage Component for Alignment Controller Verification
//
// -----------------------------------------------------------------------------
// OVERVIEW:
// The `algn_coverage` class is a UVM component responsible for collecting 
// functional coverage related to the packet-splitting behavior of the 
// Alignment Controller DUT. It monitors the `algn_split_info` transactions
// generated by the reference model and records how well different combinations 
// of control and metadata parameters are exercised.
//
// -----------------------------------------------------------------------------
// FUNCTIONAL FLOW:
// 1. The reference model sends alignment split information through its analysis
//    port (of type `algn_split_info`).
// 2. The `algn_coverage` component receives this data through its analysis 
//    implementation port (`port_in_split_info`).
// 3. For each received transaction, the `write_in_split_info()` method is called.
// 4. Inside this method, the `cover_split` covergroup samples the received data.
// 5. Coverage points track key parameters such as control offset, control size,
//    metadata offset, metadata size, and number of bytes required.
// 6. A cross coverage (`all`) captures valid combinations of these fields.
// 7. Optional debug functionality prints coverage percentages at the end of 
//    simulation (in `report_phase`), though this should not be used in 
//    production-level environments.
//
// -----------------------------------------------------------------------------
// STRUCTURE:
//  - Analysis port: `port_in_split_info`
//  - Covergroup: `cover_split`
//  - Methods:
//       * new()                : Constructor, creates covergroup and ports.
//       * write_in_split_info(): Samples the covergroup on each transaction.
//       * handle_reset()       : Placeholder for reset-related coverage logic.
//       * coverage2string()    : Formats coverage results as a string (debug only).
//       * report_phase()       : Prints coverage summary at simulation end.
//
// -----------------------------------------------------------------------------
// NOTES:
//  - This component implements `uvm_ext_reset_handler_if` to integrate 
//    with environments that broadcast resets to components.
//  - Coverage values printed in `report_phase()` are only for quick visualization 
//    and debugging (not suitable for real regressions).
///////////////////////////////////////////////////////////////////////////////

`ifndef ALGN_COVERAGE_SV
`define ALGN_COVERAGE_SV

  // Declare an analysis implementation for receiving split information
  `uvm_analysis_imp_decl(_in_split_info)

  class algn_coverage extends uvm_component implements uvm_ext_reset_handler_if;

    //--------------------------------------------------------------------------
    // Analysis implementation port
    //--------------------------------------------------------------------------
    // Used to receive split information (algn_split_info) from the model.
    // Each received transaction triggers a call to write_in_split_info().
    uvm_analysis_imp_in_split_info#(algn_split_info, algn_coverage) port_in_split_info;

    //--------------------------------------------------------------------------
    // Covergroup: cover_split
    //--------------------------------------------------------------------------
    // Tracks functional coverage of key fields in algn_split_info and
    // their combinations.
    covergroup cover_split with function sample(algn_split_info info);
      option.per_instance = 1; // Unique instance per component

      // Coverpoint: CTRL offset value
      ctrl_offset : coverpoint info.ctrl_offset {
        option.comment = "Value of CTRL.OFFSET";
        bins values[] = {[0:3]};
      }

      // Coverpoint: CTRL size value
      ctrl_size : coverpoint info.ctrl_size {
        option.comment = "Value of CTRL.SIZE";
        bins values[] = {[1:4]};
      }

      // Coverpoint: MD transaction offset
      md_offset : coverpoint info.md_offset {
        option.comment = "Value of the MD transaction offset";
        bins values[] = {[0:3]};
      }

      // Coverpoint: MD transaction size
      md_size : coverpoint info.md_size {
        option.comment = "Value of the MD transaction size";
        bins values[] = {[1:4]};
      }

      // Coverpoint: Number of bytes needed during the split
      num_bytes_needed : coverpoint info.num_bytes_needed {
        option.comment = "Number of bytes needed during the split";
        bins values[] = {[1:3]};
      }

      // Cross coverage: Valid combinations of all parameters
      all : cross ctrl_offset, ctrl_size, md_offset, md_size, num_bytes_needed {
        // Ignore illegal or invalid combinations from coverage
        ignore_bins ignore_ctrl = 
          (binsof(ctrl_offset) intersect {0} && binsof(ctrl_size) intersect {3})       ||
          (binsof(ctrl_offset) intersect {1} && binsof(ctrl_size) intersect {2, 3, 4}) ||
          (binsof(ctrl_offset) intersect {2} && binsof(ctrl_size) intersect {3, 4})    ||
          (binsof(ctrl_offset) intersect {3} && binsof(ctrl_size) intersect {2, 3, 4});
        // TODO: Add additional invalid combinations as required.
      }

    endgroup : cover_split

    //--------------------------------------------------------------------------
    // Factory registration
    //--------------------------------------------------------------------------
    `uvm_component_utils(algn_coverage)

    //--------------------------------------------------------------------------
    // Constructor
    //--------------------------------------------------------------------------
    function new(string name = "", uvm_component parent);
      super.new(name, parent);

      // Create analysis implementation port
      port_in_split_info = new("port_in_split_info", this);

      // Create and name the covergroup instance
      cover_split = new();
      cover_split.set_inst_name($sformatf("%0s_%0s", get_full_name(), "cover_split"));
    endfunction : new

    //--------------------------------------------------------------------------
    // write_in_split_info()
    //--------------------------------------------------------------------------
    // Triggered automatically when split info is received via analysis port.
    // Samples the covergroup with the received algn_split_info data.
    virtual function void write_in_split_info(algn_split_info info);
      cover_split.sample(info);
    endfunction : write_in_split_info

    //--------------------------------------------------------------------------
    // handle_reset()
    //--------------------------------------------------------------------------
    // Placeholder for handling reset events. Can be extended to clear 
    // internal data or reset coverage collection if required.
    virtual function void handle_reset(uvm_phase phase);
      // No operation for now.
    endfunction : handle_reset

    //--------------------------------------------------------------------------
    // coverage2string()
    //--------------------------------------------------------------------------
    // Utility function to convert coverage metrics into formatted string output.
    // Used only for quick debug visualization in simulation logs.
    virtual function string coverage2string();
      string result = {
        $sformatf("\n   cover_split:            %03.2f%%", cover_split.get_inst_coverage()),
        $sformatf("\n      ctrl_offset:         %03.2f%%", cover_split.ctrl_offset.get_inst_coverage()),
        $sformatf("\n      ctrl_size:           %03.2f%%", cover_split.ctrl_size.get_inst_coverage()),
        $sformatf("\n      md_offset:           %03.2f%%", cover_split.md_offset.get_inst_coverage()),
        $sformatf("\n      md_size:             %03.2f%%", cover_split.md_size.get_inst_coverage()),
        $sformatf("\n      num_bytes_needed:    %03.2f%%", cover_split.num_bytes_needed.get_inst_coverage()),
        $sformatf("\n      all:                 %03.2f%%", cover_split.all.get_inst_coverage())
      };
      return result;
    endfunction : coverage2string

    //--------------------------------------------------------------------------
    // report_phase()
    //--------------------------------------------------------------------------
    // Prints summary coverage results at the end of the simulation.
    // NOTE: For demonstration/debug only; not suitable for production use.
    virtual function void report_phase(uvm_phase phase);

      // Print coverage summary
      `uvm_info("COVERAGE", $sformatf("\nCoverage: %0s", coverage2string()), UVM_DEBUG)

      super.report_phase(phase);
    endfunction : report_phase

  endclass : algn_coverage

`endif
