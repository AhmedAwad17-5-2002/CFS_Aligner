///////////////////////////////////////////////////////////////////////////////
// File:        algn_virtual_sequence_slow_pace.sv
// Author:      Ahmed Awad-Allah Mohamed
// Date:        12/10/2025
// Description: 
// -----------------------------------------------------------------------------
// UVM Virtual Sequence: algn_virtual_sequence_slow_pace
// -----------------------------------------------------------------------------
// PURPOSE & FLOW:
// This virtual sequence coordinates and controls both RX and TX sequences of
// the Alignment Controller verification environment under a *slow-paced* 
// operation mode.
//
// It is designed to:
//  - Stimulate the DUT’s RX interface (via md_master_simple_sequence) with 
//    controlled MD packet data based on alignment width and register 
//    configuration.
//  - Monitor and validate TX responses (via md_slave_simple_sequence) that 
//    reflect the aligned output generated by the DUT.
//
// FLOW OVERVIEW:
//  1. Retrieve the alignment configuration values from the model and register
//     block (ALGN_DATA_WIDTH, CTRL.SIZE).
//  2. Launch the RX and TX sequences *concurrently* using a `fork...join`
//     block, allowing data push and response check to overlap.
//  3. On RX side:
//       - Generate MD packets whose data sizes and offsets are constrained
//         based on DUT configuration (ensuring valid packet boundaries).
//  4. On TX side:
//       - Consume pending RX items.
//       - Calculate how many TX items are expected per RX transfer.
//       - Generate TX responses with proper result signaling:
//           • MD_OKAY for valid aligned chunks.
//           • MD_ERR on the last chunk if the DUT signals an error.
//
// The “slow pace” term indicates that transactions are spaced or controlled to
// avoid high-throughput bursts—useful for debugging timing-sensitive alignment
// behavior.
//
// This sequence is built on top of the base virtual sequence 
// `algn_virtual_sequence_base`, inheriting common handles and configuration 
// access paths (e.g., `p_sequencer.my_algn_model`).
///////////////////////////////////////////////////////////////////////////////

`ifndef ALGN_VIRTUAL_SEQUENCE_SLOW_PACE_SV
`define ALGN_VIRTUAL_SEQUENCE_SLOW_PACE_SV

//------------------------------------------------------------------------------
// Class: algn_virtual_sequence_slow_pace
//------------------------------------------------------------------------------
// Extends: algn_virtual_sequence_base
// Implements a virtual sequence controlling both RX and TX sides
// of the DUT for the slow-paced alignment scenario.
//------------------------------------------------------------------------------
class algn_virtual_sequence_slow_pace extends algn_virtual_sequence_base;

  // Register with UVM factory to allow creation using type_id::create()
  `uvm_object_utils(algn_virtual_sequence_slow_pace)

  //--------------------------------------------------------------------------
  // Constructor
  //--------------------------------------------------------------------------
  function new(string name = "");
    super.new(name);
  endfunction

  //--------------------------------------------------------------------------
  // Task: body
  //--------------------------------------------------------------------------
  // - Main virtual sequence execution.
  // - Launches RX and TX stimulus concurrently.
  // - Controls data constraints and expected DUT responses.
  //--------------------------------------------------------------------------
  virtual task body();

    md_master_simple_sequence rx_sequence; // RX (Master) sequence handle

    fork
      //----------------------------------------------------------------------
      // RX Sequence Thread
      //----------------------------------------------------------------------
      begin
        // Retrieve configuration values from model and register block
        int unsigned algn_data_width = p_sequencer.my_algn_model.my_model_config.get_algn_data_width();
        int unsigned ctrl_size       = p_sequencer.my_algn_model.my_reg_block.CTRL.SIZE.get_mirrored_value();

        // Drive RX side with constrained data packet
        // Constraints ensure:
        //  1. Data is aligned with algn_data_width
        //  2. Size and offset are within legal bounds
        //  3. Data is large enough relative to CTRL.SIZE
        `uvm_do_on_with(rx_sequence, p_sequencer.md_rx_sequencer, {
          ((algn_data_width / 8) + my_md_drv_master_item.offset) % my_md_drv_master_item.data.size() == 0;
          (my_md_drv_master_item.data.size() + my_md_drv_master_item.offset) <= (algn_data_width / 8);
          my_md_drv_master_item.data.size() >= ctrl_size;
        })
      end

      //----------------------------------------------------------------------
      // TX Sequence Thread
      //----------------------------------------------------------------------
      begin
        int unsigned tx_item_idx = 0;
        int unsigned num_tx_items;

        do begin
          md_slave_simple_sequence tx_sequence;  // TX (Slave) sequence handle
          md_mon_item item_mon;                  // Monitored item from TX FIFO

          // Wait and fetch a pending item monitored from RX side
          p_sequencer.md_tx_sequencer.pending_items.get(item_mon);

          // Compute number of expected TX items per RX data block
          num_tx_items = rx_sequence.my_md_drv_master_item.data.size() /
                         p_sequencer.my_algn_model.my_reg_block.CTRL.SIZE.get_mirrored_value();

          // Drive TX sequence with response logic:
          // - For single item: MD_OKAY
          // - For multiple items: OKAY for all but last, which returns MD_ERR
          `uvm_do_on_with(tx_sequence, p_sequencer.md_tx_sequencer, {
            num_tx_items == 1                                     -> my_md_drv_slave_item.response == MD_OKAY;
            num_tx_items > 1 && tx_item_idx <  (num_tx_items - 1) -> my_md_drv_slave_item.response == MD_OKAY;
            num_tx_items > 1 && tx_item_idx == (num_tx_items - 1) -> my_md_drv_slave_item.response == MD_ERR;
          })

          tx_item_idx++;
        end while(tx_item_idx < num_tx_items);
      end
    join  // Synchronize RX and TX threads

  endtask : body

endclass : algn_virtual_sequence_slow_pace

`endif
